digraph {
	<__main__.Node object at 0x00000168B5CFA7F0> [label=outlook]
	<__main__.Node object at 0x00000168B5CFA278> [label=humidity]
	<__main__.Node object at 0x00000168B5CFA7F0> -> <__main__.Node object at 0x00000168B5CFA278> [label=sunny]
	<__main__.Node object at 0x00000168B5CFA828> [label=Death]
	<__main__.Node object at 0x00000168B5CFA278> -> <__main__.Node object at 0x00000168B5CFA828> [label=high]
	<__main__.Node object at 0x00000168B5CFA6A0> [label=Survived]
	<__main__.Node object at 0x00000168B5CFA278> -> <__main__.Node object at 0x00000168B5CFA6A0> [label=normal]
	<__main__.Node object at 0x00000168B5C91208> [label=Survived]
	<__main__.Node object at 0x00000168B5CFA7F0> -> <__main__.Node object at 0x00000168B5C91208> [label=overcast]
	<__main__.Node object at 0x00000168B5CFA748> [label=wind]
	<__main__.Node object at 0x00000168B5CFA7F0> -> <__main__.Node object at 0x00000168B5CFA748> [label=rain]
	<__main__.Node object at 0x00000168B5CFA438> [label=Survived]
	<__main__.Node object at 0x00000168B5CFA748> -> <__main__.Node object at 0x00000168B5CFA438> [label=weak]
	<__main__.Node object at 0x00000168B5CFAA20> [label=Death]
	<__main__.Node object at 0x00000168B5CFA748> -> <__main__.Node object at 0x00000168B5CFAA20> [label=strong]
}
