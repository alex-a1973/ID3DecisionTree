digraph {
	<__main__.Node object at 0x00000215829AEDA0> [label=Sex]
	<__main__.Node object at 0x00000215829ACA90> [label=Age]
	<__main__.Node object at 0x00000215829AEDA0> -> <__main__.Node object at 0x00000215829ACA90> [label=male]
	<__main__.Node object at 0x00000215829AC160> [label=Pclass]
	<__main__.Node object at 0x00000215829ACA90> -> <__main__.Node object at 0x00000215829AC160> [label=adults]
	<__main__.Node object at 0x00000215829AC470> [label=Embarked]
	<__main__.Node object at 0x00000215829AC160> -> <__main__.Node object at 0x00000215829AC470> [label=3]
	<__main__.Node object at 0x00000215839A97F0> [label=Fare]
	<__main__.Node object at 0x00000215829AC470> -> <__main__.Node object at 0x00000215839A97F0> [label=Q]
	<__main__.Node object at 0x00000215829ACA58> [label=Death]
	<__main__.Node object at 0x00000215839A97F0> -> <__main__.Node object at 0x00000215829ACA58> [label="middle class"]
	<__main__.Node object at 0x00000215829AE198> [label=SibSp]
	<__main__.Node object at 0x00000215839A97F0> -> <__main__.Node object at 0x00000215829AE198> [label=poor]
	<__main__.Node object at 0x00000215829AE0F0> [label=Death]
	<__main__.Node object at 0x00000215829AE198> -> <__main__.Node object at 0x00000215829AE0F0> [label=1]
	<__main__.Node object at 0x00000215829AE1D0> [label=Parch]
	<__main__.Node object at 0x00000215829AE198> -> <__main__.Node object at 0x00000215829AE1D0> [label=0]
	<__main__.Node object at 0x00000215839A9630> [label=Death]
	<__main__.Node object at 0x00000215829AE1D0> -> <__main__.Node object at 0x00000215839A9630> [label=0]
	<__main__.Node object at 0x00000215829AC0B8> [label=Fare]
	<__main__.Node object at 0x00000215829AC470> -> <__main__.Node object at 0x00000215829AC0B8> [label=S]
	<__main__.Node object at 0x00000215839A9358> [label=SibSp]
	<__main__.Node object at 0x00000215829AC0B8> -> <__main__.Node object at 0x00000215839A9358> [label=poor]
	<__main__.Node object at 0x00000215839A9BA8> [label=Parch]
	<__main__.Node object at 0x00000215839A9358> -> <__main__.Node object at 0x00000215839A9BA8> [label=0]
	<__main__.Node object at 0x00000215839A91D0> [label=Death]
	<__main__.Node object at 0x00000215839A9BA8> -> <__main__.Node object at 0x00000215839A91D0> [label=0]
	<__main__.Node object at 0x00000215839A9A90> [label=Death]
	<__main__.Node object at 0x00000215839A9BA8> -> <__main__.Node object at 0x00000215839A9A90> [label=1]
	<__main__.Node object at 0x00000215839A9B00> [label=Parch]
	<__main__.Node object at 0x00000215839A9358> -> <__main__.Node object at 0x00000215839A9B00> [label=1]
	<__main__.Node object at 0x00000215839A94A8> [label=Death]
	<__main__.Node object at 0x00000215839A9B00> -> <__main__.Node object at 0x00000215839A94A8> [label=0]
	<__main__.Node object at 0x00000215839A92B0> [label=Death]
	<__main__.Node object at 0x00000215839A9358> -> <__main__.Node object at 0x00000215839A92B0> [label=2]
	<__main__.Node object at 0x00000215839A95C0> [label=Death]
	<__main__.Node object at 0x00000215829AC0B8> -> <__main__.Node object at 0x00000215839A95C0> [label="middle class"]
	<__main__.Node object at 0x00000215839A9898> [label=SibSp]
	<__main__.Node object at 0x00000215829AC0B8> -> <__main__.Node object at 0x00000215839A9898> [label="upper class"]
	<__main__.Node object at 0x00000215839A9AC8> [label=Death]
	<__main__.Node object at 0x00000215839A9898> -> <__main__.Node object at 0x00000215839A9AC8> [label=8]
	<__main__.Node object at 0x00000215839A9B38> [label=Parch]
	<__main__.Node object at 0x00000215839A9898> -> <__main__.Node object at 0x00000215839A9B38> [label=0]
	<__main__.Node object at 0x00000215839A90B8> [label=Survived]
	<__main__.Node object at 0x00000215839A9B38> -> <__main__.Node object at 0x00000215839A90B8> [label=0]
	<__main__.Node object at 0x00000215829AE588> [label=Parch]
	<__main__.Node object at 0x00000215829AC470> -> <__main__.Node object at 0x00000215829AE588> [label=C]
	<__main__.Node object at 0x00000215829ACB00> [label=SibSp]
	<__main__.Node object at 0x00000215829AE588> -> <__main__.Node object at 0x00000215829ACB00> [label=0]
	<__main__.Node object at 0x00000215839A9940> [label=Fare]
	<__main__.Node object at 0x00000215829ACB00> -> <__main__.Node object at 0x00000215839A9940> [label=0]
	<__main__.Node object at 0x0000021582964C18> [label=Death]
	<__main__.Node object at 0x00000215839A9940> -> <__main__.Node object at 0x0000021582964C18> [label=poor]
	<__main__.Node object at 0x0000021582964BE0> [label=Survived]
	<__main__.Node object at 0x00000215839A9940> -> <__main__.Node object at 0x0000021582964BE0> [label="middle class"]
	<__main__.Node object at 0x00000215839A9860> [label=Death]
	<__main__.Node object at 0x00000215829ACB00> -> <__main__.Node object at 0x00000215839A9860> [label=2]
	<__main__.Node object at 0x00000215839A99E8> [label=Death]
	<__main__.Node object at 0x00000215829ACB00> -> <__main__.Node object at 0x00000215839A99E8> [label=1]
	<__main__.Node object at 0x00000215839A92E8> [label=Survived]
	<__main__.Node object at 0x00000215829AE588> -> <__main__.Node object at 0x00000215839A92E8> [label=1]
	<__main__.Node object at 0x00000215829AC4E0> [label=SibSp]
	<__main__.Node object at 0x00000215829AC160> -> <__main__.Node object at 0x00000215829AC4E0> [label=2]
	<__main__.Node object at 0x00000215839A9748> [label=Fare]
	<__main__.Node object at 0x00000215829AC4E0> -> <__main__.Node object at 0x00000215839A9748> [label=0]
	<__main__.Node object at 0x00000215839A9DD8> [label=Embarked]
	<__main__.Node object at 0x00000215839A9748> -> <__main__.Node object at 0x00000215839A9DD8> [label="middle class"]
	<__main__.Node object at 0x0000021582964668> [label=Parch]
	<__main__.Node object at 0x00000215839A9DD8> -> <__main__.Node object at 0x0000021582964668> [label=S]
	<__main__.Node object at 0x0000021582964DD8> [label=Death]
	<__main__.Node object at 0x0000021582964668> -> <__main__.Node object at 0x0000021582964DD8> [label=0]
	<__main__.Node object at 0x0000021582964B38> [label=Death]
	<__main__.Node object at 0x0000021582964668> -> <__main__.Node object at 0x0000021582964B38> [label=2]
	<__main__.Node object at 0x00000215829640F0> [label=Death]
	<__main__.Node object at 0x0000021582964668> -> <__main__.Node object at 0x00000215829640F0> [label=1]
	<__main__.Node object at 0x0000021582964860> [label=Death]
	<__main__.Node object at 0x00000215839A9DD8> -> <__main__.Node object at 0x0000021582964860> [label=Q]
	<__main__.Node object at 0x0000021582964240> [label=Death]
	<__main__.Node object at 0x00000215839A9DD8> -> <__main__.Node object at 0x0000021582964240> [label=C]
	<__main__.Node object at 0x00000215839A9400> [label=Death]
	<__main__.Node object at 0x00000215839A9748> -> <__main__.Node object at 0x00000215839A9400> [label="upper class"]
	<__main__.Node object at 0x00000215839A9160> [label=Death]
	<__main__.Node object at 0x00000215839A9748> -> <__main__.Node object at 0x00000215839A9160> [label=poor]
	<__main__.Node object at 0x00000215839A9390> [label=Death]
	<__main__.Node object at 0x00000215829AC4E0> -> <__main__.Node object at 0x00000215839A9390> [label=1]
	<__main__.Node object at 0x00000215839A9048> [label=Death]
	<__main__.Node object at 0x00000215829AC4E0> -> <__main__.Node object at 0x00000215839A9048> [label=2]
	<__main__.Node object at 0x00000215829ACAC8> [label=SibSp]
	<__main__.Node object at 0x00000215829AC160> -> <__main__.Node object at 0x00000215829ACAC8> [label=1]
	<__main__.Node object at 0x00000215839A96D8> [label=Fare]
	<__main__.Node object at 0x00000215829ACAC8> -> <__main__.Node object at 0x00000215839A96D8> [label=0]
	<__main__.Node object at 0x00000215839A9A58> [label=Parch]
	<__main__.Node object at 0x00000215839A96D8> -> <__main__.Node object at 0x00000215839A9A58> [label="middle class"]
	<__main__.Node object at 0x0000021582964748> [label=Embarked]
	<__main__.Node object at 0x00000215839A9A58> -> <__main__.Node object at 0x0000021582964748> [label=0]
	<__main__.Node object at 0x00000215829645F8> [label=Death]
	<__main__.Node object at 0x0000021582964748> -> <__main__.Node object at 0x00000215829645F8> [label=C]
	<__main__.Node object at 0x0000021582964908> [label=Death]
	<__main__.Node object at 0x0000021582964748> -> <__main__.Node object at 0x0000021582964908> [label=S]
	<__main__.Node object at 0x0000021582964518> [label=Death]
	<__main__.Node object at 0x00000215839A9A58> -> <__main__.Node object at 0x0000021582964518> [label=1]
	<__main__.Node object at 0x00000215829647F0> [label=Embarked]
	<__main__.Node object at 0x00000215839A96D8> -> <__main__.Node object at 0x00000215829647F0> [label="upper class"]
	<__main__.Node object at 0x0000021582964A90> [label=Death]
	<__main__.Node object at 0x00000215829647F0> -> <__main__.Node object at 0x0000021582964A90> [label=S]
	<__main__.Node object at 0x0000021582964470> [label=Parch]
	<__main__.Node object at 0x00000215829647F0> -> <__main__.Node object at 0x0000021582964470> [label=C]
	<__main__.Node object at 0x00000215829649E8> [label=Death]
	<__main__.Node object at 0x0000021582964470> -> <__main__.Node object at 0x00000215829649E8> [label=0]
	<__main__.Node object at 0x0000021582964390> [label=Death]
	<__main__.Node object at 0x0000021582964470> -> <__main__.Node object at 0x0000021582964390> [label=1]
	<__main__.Node object at 0x00000215829645C0> [label=Death]
	<__main__.Node object at 0x0000021582964470> -> <__main__.Node object at 0x00000215829645C0> [label=2]
	<__main__.Node object at 0x0000021582964400> [label=Death]
	<__main__.Node object at 0x00000215839A96D8> -> <__main__.Node object at 0x0000021582964400> [label=poor]
	<__main__.Node object at 0x00000215839A9278> [label=Parch]
	<__main__.Node object at 0x00000215829ACAC8> -> <__main__.Node object at 0x00000215839A9278> [label=1]
	<__main__.Node object at 0x00000215839A99B0> [label=Embarked]
	<__main__.Node object at 0x00000215839A9278> -> <__main__.Node object at 0x00000215839A99B0> [label=0]
	<__main__.Node object at 0x00000215839F15C0> [label=Fare]
	<__main__.Node object at 0x00000215839A99B0> -> <__main__.Node object at 0x00000215839F15C0> [label=S]
	<__main__.Node object at 0x00000215839F14E0> [label=Death]
	<__main__.Node object at 0x00000215839F15C0> -> <__main__.Node object at 0x00000215839F14E0> [label="upper class"]
	<__main__.Node object at 0x00000215839F1080> [label=Fare]
	<__main__.Node object at 0x00000215839A99B0> -> <__main__.Node object at 0x00000215839F1080> [label=C]
	<__main__.Node object at 0x00000215839F1048> [label=Survived]
	<__main__.Node object at 0x00000215839F1080> -> <__main__.Node object at 0x00000215839F1048> [label="upper class"]
	<__main__.Node object at 0x0000021582964D30> [label=Death]
	<__main__.Node object at 0x00000215839A9278> -> <__main__.Node object at 0x0000021582964D30> [label=4]
	<__main__.Node object at 0x0000021582964828> [label=Embarked]
	<__main__.Node object at 0x00000215839A9278> -> <__main__.Node object at 0x0000021582964828> [label=1]
	<__main__.Node object at 0x00000215839F1588> [label=Fare]
	<__main__.Node object at 0x0000021582964828> -> <__main__.Node object at 0x00000215839F1588> [label=C]
	<__main__.Node object at 0x00000215839F1438> [label=Survived]
	<__main__.Node object at 0x00000215839F1588> -> <__main__.Node object at 0x00000215839F1438> [label="upper class"]
	<__main__.Node object at 0x00000215839F10B8> [label=Survived]
	<__main__.Node object at 0x0000021582964828> -> <__main__.Node object at 0x00000215839F10B8> [label=S]
	<__main__.Node object at 0x00000215829643C8> [label=Survived]
	<__main__.Node object at 0x00000215839A9278> -> <__main__.Node object at 0x00000215829643C8> [label=2]
	<__main__.Node object at 0x00000215839A97B8> [label=Death]
	<__main__.Node object at 0x00000215829ACAC8> -> <__main__.Node object at 0x00000215839A97B8> [label=3]
	<__main__.Node object at 0x00000215839A98D0> [label=Embarked]
	<__main__.Node object at 0x00000215829ACAC8> -> <__main__.Node object at 0x00000215839A98D0> [label=2]
	<__main__.Node object at 0x0000021582964CF8> [label=Death]
	<__main__.Node object at 0x00000215839A98D0> -> <__main__.Node object at 0x0000021582964CF8> [label=Q]
	<__main__.Node object at 0x0000021582964898> [label=Survived]
	<__main__.Node object at 0x00000215839A98D0> -> <__main__.Node object at 0x0000021582964898> [label=S]
	<__main__.Node object at 0x00000215829AC0F0> [label=Parch]
	<__main__.Node object at 0x00000215829ACA90> -> <__main__.Node object at 0x00000215829AC0F0> [label=teen]
	<__main__.Node object at 0x00000215829AC8D0> [label=Death]
	<__main__.Node object at 0x00000215829AC0F0> -> <__main__.Node object at 0x00000215829AC8D0> [label=1]
	<__main__.Node object at 0x00000215829AC080> [label=Fare]
	<__main__.Node object at 0x00000215829AC0F0> -> <__main__.Node object at 0x00000215829AC080> [label=0]
	<__main__.Node object at 0x00000215839A93C8> [label=SibSp]
	<__main__.Node object at 0x00000215829AC080> -> <__main__.Node object at 0x00000215839A93C8> [label=poor]
	<__main__.Node object at 0x00000215839F1550> [label=Pclass]
	<__main__.Node object at 0x00000215839A93C8> -> <__main__.Node object at 0x00000215839F1550> [label=0]
	<__main__.Node object at 0x00000215839F15F8> [label=Embarked]
	<__main__.Node object at 0x00000215839F1550> -> <__main__.Node object at 0x00000215839F15F8> [label=3]
	<__main__.Node object at 0x00000215839F1B00> [label=Death]
	<__main__.Node object at 0x00000215839F15F8> -> <__main__.Node object at 0x00000215839F1B00> [label=S]
	<__main__.Node object at 0x00000215839F1358> [label=Death]
	<__main__.Node object at 0x00000215839A93C8> -> <__main__.Node object at 0x00000215839F1358> [label=1]
	<__main__.Node object at 0x0000021582964588> [label=Death]
	<__main__.Node object at 0x00000215829AC080> -> <__main__.Node object at 0x0000021582964588> [label="upper class"]
	<__main__.Node object at 0x0000021582964198> [label=Death]
	<__main__.Node object at 0x00000215829AC080> -> <__main__.Node object at 0x0000021582964198> [label="middle class"]
	<__main__.Node object at 0x00000215839A9550> [label=Death]
	<__main__.Node object at 0x00000215829AC0F0> -> <__main__.Node object at 0x00000215839A9550> [label=3]
	<__main__.Node object at 0x00000215829AC048> [label=Pclass]
	<__main__.Node object at 0x00000215829AC0F0> -> <__main__.Node object at 0x00000215829AC048> [label=2]
	<__main__.Node object at 0x00000215839F12B0> [label=Survived]
	<__main__.Node object at 0x00000215829AC048> -> <__main__.Node object at 0x00000215839F12B0> [label=1]
	<__main__.Node object at 0x00000215839F14A8> [label=Death]
	<__main__.Node object at 0x00000215829AC048> -> <__main__.Node object at 0x00000215839F14A8> [label=3]
	<__main__.Node object at 0x0000021582964320> [label=SibSp]
	<__main__.Node object at 0x00000215829ACA90> -> <__main__.Node object at 0x0000021582964320> [label=child]
	<__main__.Node object at 0x00000215829647B8> [label=Parch]
	<__main__.Node object at 0x0000021582964320> -> <__main__.Node object at 0x00000215829647B8> [label=4]
	<__main__.Node object at 0x00000215839A9438> [label=Death]
	<__main__.Node object at 0x00000215829647B8> -> <__main__.Node object at 0x00000215839A9438> [label=1]
	<__main__.Node object at 0x00000215839F1320> [label=Pclass]
	<__main__.Node object at 0x00000215829647B8> -> <__main__.Node object at 0x00000215839F1320> [label=2]
	<__main__.Node object at 0x00000215839F1710> [label=Fare]
	<__main__.Node object at 0x00000215839F1320> -> <__main__.Node object at 0x00000215839F1710> [label=3]
	<__main__.Node object at 0x00000215839F1E48> [label=Embarked]
	<__main__.Node object at 0x00000215839F1710> -> <__main__.Node object at 0x00000215839F1E48> [label="middle class"]
	<__main__.Node object at 0x00000215839F1FD0> [label=Death]
	<__main__.Node object at 0x00000215839F1E48> -> <__main__.Node object at 0x00000215839F1FD0> [label=S]
	<__main__.Node object at 0x00000215829ACE80> [label=Survived]
	<__main__.Node object at 0x0000021582964320> -> <__main__.Node object at 0x00000215829ACE80> [label=2]
	<__main__.Node object at 0x00000215839F1278> [label=Survived]
	<__main__.Node object at 0x0000021582964320> -> <__main__.Node object at 0x00000215839F1278> [label=1]
	<__main__.Node object at 0x00000215839F1828> [label=Death]
	<__main__.Node object at 0x0000021582964320> -> <__main__.Node object at 0x00000215839F1828> [label=3]
	<__main__.Node object at 0x00000215839F17B8> [label=Parch]
	<__main__.Node object at 0x0000021582964320> -> <__main__.Node object at 0x00000215839F17B8> [label=0]
	<__main__.Node object at 0x00000215839F1BE0> [label=Death]
	<__main__.Node object at 0x00000215839F17B8> -> <__main__.Node object at 0x00000215839F1BE0> [label=0]
	<__main__.Node object at 0x00000215839F1898> [label=Survived]
	<__main__.Node object at 0x00000215839F17B8> -> <__main__.Node object at 0x00000215839F1898> [label=1]
	<__main__.Node object at 0x00000215839F1C18> [label=Survived]
	<__main__.Node object at 0x00000215839F17B8> -> <__main__.Node object at 0x00000215839F1C18> [label=2]
	<__main__.Node object at 0x00000215839F1AC8> [label=Death]
	<__main__.Node object at 0x0000021582964320> -> <__main__.Node object at 0x00000215839F1AC8> [label=5]
	<__main__.Node object at 0x00000215829ACC50> [label=Fare]
	<__main__.Node object at 0x00000215829ACA90> -> <__main__.Node object at 0x00000215829ACC50> [label=elderly]
	<__main__.Node object at 0x00000215839F16A0> [label=Pclass]
	<__main__.Node object at 0x00000215829ACC50> -> <__main__.Node object at 0x00000215839F16A0> [label="middle class"]
	<__main__.Node object at 0x00000215839F1160> [label=Death]
	<__main__.Node object at 0x00000215839F16A0> -> <__main__.Node object at 0x00000215839F1160> [label=2]
	<__main__.Node object at 0x00000215839F19E8> [label=Embarked]
	<__main__.Node object at 0x00000215839F16A0> -> <__main__.Node object at 0x00000215839F19E8> [label=1]
	<__main__.Node object at 0x00000215839F1128> [label=SibSp]
	<__main__.Node object at 0x00000215839F19E8> -> <__main__.Node object at 0x00000215839F1128> [label=S]
	<__main__.Node object at 0x00000215829640B8> [label=Parch]
	<__main__.Node object at 0x00000215839F1128> -> <__main__.Node object at 0x00000215829640B8> [label=0]
	<__main__.Node object at 0x00000215839A9978> [label=Survived]
	<__main__.Node object at 0x00000215829640B8> -> <__main__.Node object at 0x00000215839A9978> [label=0]
	<__main__.Node object at 0x00000215839F1198> [label=Death]
	<__main__.Node object at 0x00000215839F19E8> -> <__main__.Node object at 0x00000215839F1198> [label=C]
	<__main__.Node object at 0x00000215839F1630> [label=Death]
	<__main__.Node object at 0x00000215829ACC50> -> <__main__.Node object at 0x00000215839F1630> [label=poor]
	<__main__.Node object at 0x00000215839F10F0> [label=Death]
	<__main__.Node object at 0x00000215829ACC50> -> <__main__.Node object at 0x00000215839F10F0> [label="upper class"]
	<__main__.Node object at 0x00000215829AC5F8> [label=Pclass]
	<__main__.Node object at 0x00000215829AEDA0> -> <__main__.Node object at 0x00000215829AC5F8> [label=female]
	<__main__.Node object at 0x00000215829AC3C8> [label=Parch]
	<__main__.Node object at 0x00000215829AC5F8> -> <__main__.Node object at 0x00000215829AC3C8> [label=3]
	<__main__.Node object at 0x00000215839F1F28> [label=Embarked]
	<__main__.Node object at 0x00000215829AC3C8> -> <__main__.Node object at 0x00000215839F1F28> [label=0]
	<__main__.Node object at 0x00000215839F1CC0> [label=SibSp]
	<__main__.Node object at 0x00000215839F1F28> -> <__main__.Node object at 0x00000215839F1CC0> [label=S]
	<__main__.Node object at 0x00000215839A9710> [label=Fare]
	<__main__.Node object at 0x00000215839F1CC0> -> <__main__.Node object at 0x00000215839A9710> [label=0]
	<__main__.Node object at 0x00000215839A94E0> [label=Age]
	<__main__.Node object at 0x00000215839A9710> -> <__main__.Node object at 0x00000215839A94E0> [label=poor]
	<__main__.Node object at 0x00000215839EA160> [label=Death]
	<__main__.Node object at 0x00000215839A94E0> -> <__main__.Node object at 0x00000215839EA160> [label=adults]
	<__main__.Node object at 0x00000215839EA128> [label=Survived]
	<__main__.Node object at 0x00000215839A94E0> -> <__main__.Node object at 0x00000215839EA128> [label=teen]
	<__main__.Node object at 0x00000215839A9BE0> [label=Survived]
	<__main__.Node object at 0x00000215839A9710> -> <__main__.Node object at 0x00000215839A9BE0> [label="middle class"]
	<__main__.Node object at 0x00000215839A9080> [label=Fare]
	<__main__.Node object at 0x00000215839F1CC0> -> <__main__.Node object at 0x00000215839A9080> [label=1]
	<__main__.Node object at 0x00000215839A9668> [label=Age]
	<__main__.Node object at 0x00000215839A9080> -> <__main__.Node object at 0x00000215839A9668> [label="middle class"]
	<__main__.Node object at 0x00000215839EA240> [label=Survived]
	<__main__.Node object at 0x00000215839A9668> -> <__main__.Node object at 0x00000215839EA240> [label=adults]
	<__main__.Node object at 0x00000215839A9E10> [label=Age]
	<__main__.Node object at 0x00000215839A9080> -> <__main__.Node object at 0x00000215839A9E10> [label=poor]
	<__main__.Node object at 0x00000215839EA0F0> [label=Death]
	<__main__.Node object at 0x00000215839A9E10> -> <__main__.Node object at 0x00000215839EA0F0> [label=adults]
	<__main__.Node object at 0x0000021582943CC0> [label=Survived]
	<__main__.Node object at 0x00000215839F1CC0> -> <__main__.Node object at 0x0000021582943CC0> [label=3]
	<__main__.Node object at 0x00000215839A9198> [label=Death]
	<__main__.Node object at 0x00000215839F1CC0> -> <__main__.Node object at 0x00000215839A9198> [label=2]
	<__main__.Node object at 0x0000021582964AC8> [label=SibSp]
	<__main__.Node object at 0x00000215839F1F28> -> <__main__.Node object at 0x0000021582964AC8> [label=Q]
	<__main__.Node object at 0x00000215839A9828> [label=Survived]
	<__main__.Node object at 0x0000021582964AC8> -> <__main__.Node object at 0x00000215839A9828> [label=1]
	<__main__.Node object at 0x0000021582964080> [label=Age]
	<__main__.Node object at 0x0000021582964AC8> -> <__main__.Node object at 0x0000021582964080> [label=0]
	<__main__.Node object at 0x00000215839EA4A8> [label=Fare]
	<__main__.Node object at 0x0000021582964080> -> <__main__.Node object at 0x00000215839EA4A8> [label=adults]
	<__main__.Node object at 0x00000215839EA6D8> [label=Survived]
	<__main__.Node object at 0x00000215839EA4A8> -> <__main__.Node object at 0x00000215839EA6D8> [label=poor]
	<__main__.Node object at 0x00000215839EA320> [label=Fare]
	<__main__.Node object at 0x0000021582964080> -> <__main__.Node object at 0x00000215839EA320> [label=teen]
	<__main__.Node object at 0x00000215839EA748> [label=Survived]
	<__main__.Node object at 0x00000215839EA320> -> <__main__.Node object at 0x00000215839EA748> [label=poor]
	<__main__.Node object at 0x0000021582964B70> [label=Survived]
	<__main__.Node object at 0x0000021582964AC8> -> <__main__.Node object at 0x0000021582964B70> [label=2]
	<__main__.Node object at 0x00000215839A9518> [label=Fare]
	<__main__.Node object at 0x00000215839F1F28> -> <__main__.Node object at 0x00000215839A9518> [label=C]
	<__main__.Node object at 0x00000215829AE0B8> [label=Survived]
	<__main__.Node object at 0x00000215839A9518> -> <__main__.Node object at 0x00000215829AE0B8> [label=poor]
	<__main__.Node object at 0x00000215829AE128> [label=Age]
	<__main__.Node object at 0x00000215839A9518> -> <__main__.Node object at 0x00000215829AE128> [label="middle class"]
	<__main__.Node object at 0x00000215839EA860> [label=SibSp]
	<__main__.Node object at 0x00000215829AE128> -> <__main__.Node object at 0x00000215839EA860> [label=teen]
	<__main__.Node object at 0x00000215829AE240> [label=Survived]
	<__main__.Node object at 0x00000215839EA860> -> <__main__.Node object at 0x00000215829AE240> [label=1]
	<__main__.Node object at 0x0000021582964A20> [label=Death]
	<__main__.Node object at 0x00000215839EA860> -> <__main__.Node object at 0x0000021582964A20> [label=0]
	<__main__.Node object at 0x00000215829ACBA8> [label=Death]
	<__main__.Node object at 0x00000215829AE128> -> <__main__.Node object at 0x00000215829ACBA8> [label=adults]
	<__main__.Node object at 0x00000215829AC9B0> [label=SibSp]
	<__main__.Node object at 0x00000215829AC3C8> -> <__main__.Node object at 0x00000215829AC9B0> [label=2]
	<__main__.Node object at 0x00000215839A9A20> [label=Embarked]
	<__main__.Node object at 0x00000215829AC9B0> -> <__main__.Node object at 0x00000215839A9A20> [label=0]
	<__main__.Node object at 0x00000215839F1DA0> [label=Death]
	<__main__.Node object at 0x00000215839A9A20> -> <__main__.Node object at 0x00000215839F1DA0> [label=Q]
	<__main__.Node object at 0x00000215839F1208> [label=Survived]
	<__main__.Node object at 0x00000215839A9A20> -> <__main__.Node object at 0x00000215839F1208> [label=C]
	<__main__.Node object at 0x00000215839F1470> [label=Age]
	<__main__.Node object at 0x00000215839A9A20> -> <__main__.Node object at 0x00000215839F1470> [label=S]
	<__main__.Node object at 0x00000215839EA898> [label=Fare]
	<__main__.Node object at 0x00000215839F1470> -> <__main__.Node object at 0x00000215839EA898> [label=adults]
	<__main__.Node object at 0x00000215839EAB00> [label=Survived]
	<__main__.Node object at 0x00000215839EA898> -> <__main__.Node object at 0x00000215839EAB00> [label="middle class"]
	<__main__.Node object at 0x00000215839EA940> [label=Survived]
	<__main__.Node object at 0x00000215839F1470> -> <__main__.Node object at 0x00000215839EA940> [label=child]
	<__main__.Node object at 0x00000215839F1EF0> [label=Age]
	<__main__.Node object at 0x00000215829AC9B0> -> <__main__.Node object at 0x00000215839F1EF0> [label=4]
	<__main__.Node object at 0x00000215839F17F0> [label=Fare]
	<__main__.Node object at 0x00000215839F1EF0> -> <__main__.Node object at 0x00000215839F17F0> [label=child]
	<__main__.Node object at 0x00000215839EAA90> [label=Embarked]
	<__main__.Node object at 0x00000215839F17F0> -> <__main__.Node object at 0x00000215839EAA90> [label="middle class"]
	<__main__.Node object at 0x00000215839EA518> [label=Death]
	<__main__.Node object at 0x00000215839EAA90> -> <__main__.Node object at 0x00000215839EA518> [label=S]
	<__main__.Node object at 0x00000215839A9B70> [label=Survived]
	<__main__.Node object at 0x00000215839F1EF0> -> <__main__.Node object at 0x00000215839A9B70> [label=teen]
	<__main__.Node object at 0x00000215839F1F98> [label=Death]
	<__main__.Node object at 0x00000215829AC9B0> -> <__main__.Node object at 0x00000215839F1F98> [label=8]
	<__main__.Node object at 0x00000215839F1908> [label=Death]
	<__main__.Node object at 0x00000215829AC9B0> -> <__main__.Node object at 0x00000215839F1908> [label=2]
	<__main__.Node object at 0x00000215839F1390> [label=Death]
	<__main__.Node object at 0x00000215829AC9B0> -> <__main__.Node object at 0x00000215839F1390> [label=1]
	<__main__.Node object at 0x00000215839F1EB8> [label=Death]
	<__main__.Node object at 0x00000215829AC9B0> -> <__main__.Node object at 0x00000215839F1EB8> [label=3]
	<__main__.Node object at 0x00000215839F1F60> [label=Death]
	<__main__.Node object at 0x00000215829AC9B0> -> <__main__.Node object at 0x00000215839F1F60> [label=5]
	<__main__.Node object at 0x00000215829AC2E8> [label=SibSp]
	<__main__.Node object at 0x00000215829AC3C8> -> <__main__.Node object at 0x00000215829AC2E8> [label=1]
	<__main__.Node object at 0x0000021582964048> [label=Age]
	<__main__.Node object at 0x00000215829AC2E8> -> <__main__.Node object at 0x0000021582964048> [label=0]
	<__main__.Node object at 0x00000215839EA470> [label=Embarked]
	<__main__.Node object at 0x0000021582964048> -> <__main__.Node object at 0x00000215839EA470> [label=child]
	<__main__.Node object at 0x00000215839EA278> [label=Survived]
	<__main__.Node object at 0x00000215839EA470> -> <__main__.Node object at 0x00000215839EA278> [label=C]
	<__main__.Node object at 0x00000215839EA048> [label=Fare]
	<__main__.Node object at 0x00000215839EA470> -> <__main__.Node object at 0x00000215839EA048> [label=S]
	<__main__.Node object at 0x00000215839EACF8> [label=Survived]
	<__main__.Node object at 0x00000215839EA048> -> <__main__.Node object at 0x00000215839EACF8> [label="middle class"]
	<__main__.Node object at 0x00000215839EA780> [label=Embarked]
	<__main__.Node object at 0x0000021582964048> -> <__main__.Node object at 0x00000215839EA780> [label=adults]
	<__main__.Node object at 0x00000215839EA9E8> [label=Survived]
	<__main__.Node object at 0x00000215839EA780> -> <__main__.Node object at 0x00000215839EA9E8> [label=S]
	<__main__.Node object at 0x00000215839EA668> [label=Death]
	<__main__.Node object at 0x00000215839EA780> -> <__main__.Node object at 0x00000215839EA668> [label=C]
	<__main__.Node object at 0x00000215839EAAC8> [label=Death]
	<__main__.Node object at 0x0000021582964048> -> <__main__.Node object at 0x00000215839EAAC8> [label=teen]
	<__main__.Node object at 0x0000021582964C50> [label=Death]
	<__main__.Node object at 0x00000215829AC2E8> -> <__main__.Node object at 0x0000021582964C50> [label=3]
	<__main__.Node object at 0x00000215839EAF60> [label=Age]
	<__main__.Node object at 0x00000215829AC2E8> -> <__main__.Node object at 0x00000215839EAF60> [label=1]
	<__main__.Node object at 0x00000215839EAE80> [label=Embarked]
	<__main__.Node object at 0x00000215839EAF60> -> <__main__.Node object at 0x00000215839EAE80> [label=adults]
	<__main__.Node object at 0x00000215839EAF98> [label=Fare]
	<__main__.Node object at 0x00000215839EAE80> -> <__main__.Node object at 0x00000215839EAF98> [label=S]
	<__main__.Node object at 0x0000021583A21208> [label=Death]
	<__main__.Node object at 0x00000215839EAF98> -> <__main__.Node object at 0x0000021583A21208> [label="middle class"]
	<__main__.Node object at 0x00000215839EAE48> [label=Death]
	<__main__.Node object at 0x00000215839EAE80> -> <__main__.Node object at 0x00000215839EAE48> [label=Q]
	<__main__.Node object at 0x00000215839EABA8> [label=Survived]
	<__main__.Node object at 0x00000215839EAF60> -> <__main__.Node object at 0x00000215839EABA8> [label=child]
	<__main__.Node object at 0x00000215839EAA58> [label=Survived]
	<__main__.Node object at 0x00000215829AC2E8> -> <__main__.Node object at 0x00000215839EAA58> [label=2]
	<__main__.Node object at 0x0000021582964B00> [label=Death]
	<__main__.Node object at 0x00000215829AC3C8> -> <__main__.Node object at 0x0000021582964B00> [label=5]
	<__main__.Node object at 0x00000215839F1C50> [label=SibSp]
	<__main__.Node object at 0x00000215829AC3C8> -> <__main__.Node object at 0x00000215839F1C50> [label=3]
	<__main__.Node object at 0x00000215839EA400> [label=Death]
	<__main__.Node object at 0x00000215839F1C50> -> <__main__.Node object at 0x00000215839EA400> [label=1]
	<__main__.Node object at 0x00000215839EADA0> [label=Survived]
	<__main__.Node object at 0x00000215839F1C50> -> <__main__.Node object at 0x00000215839EADA0> [label=0]
	<__main__.Node object at 0x00000215839A9780> [label=Death]
	<__main__.Node object at 0x00000215829AC3C8> -> <__main__.Node object at 0x00000215839A9780> [label=4]
	<__main__.Node object at 0x00000215839F1A58> [label=Age]
	<__main__.Node object at 0x00000215829AC5F8> -> <__main__.Node object at 0x00000215839F1A58> [label=1]
	<__main__.Node object at 0x00000215839F1668> [label=Parch]
	<__main__.Node object at 0x00000215839F1A58> -> <__main__.Node object at 0x00000215839F1668> [label=adults]
	<__main__.Node object at 0x00000215839EAEF0> [label=Fare]
	<__main__.Node object at 0x00000215839F1668> -> <__main__.Node object at 0x00000215839EAEF0> [label=0]
	<__main__.Node object at 0x0000021583A212E8> [label=Survived]
	<__main__.Node object at 0x00000215839EAEF0> -> <__main__.Node object at 0x0000021583A212E8> [label="upper class"]
	<__main__.Node object at 0x0000021583A21240> [label=Embarked]
	<__main__.Node object at 0x00000215839EAEF0> -> <__main__.Node object at 0x0000021583A21240> [label="middle class"]
	<__main__.Node object at 0x0000021583A21400> [label=Survived]
	<__main__.Node object at 0x0000021583A21240> -> <__main__.Node object at 0x0000021583A21400> [label=S]
	<__main__.Node object at 0x0000021583A21668> [label=SibSp]
	<__main__.Node object at 0x0000021583A21240> -> <__main__.Node object at 0x0000021583A21668> [label=C]
	<__main__.Node object at 0x0000021583A21198> [label=Survived]
	<__main__.Node object at 0x0000021583A21668> -> <__main__.Node object at 0x0000021583A21198> [label=0]
	<__main__.Node object at 0x0000021583A21860> [label=Survived]
	<__main__.Node object at 0x0000021583A21668> -> <__main__.Node object at 0x0000021583A21860> [label=1]
	<__main__.Node object at 0x00000215839EA2B0> [label=SibSp]
	<__main__.Node object at 0x00000215839F1668> -> <__main__.Node object at 0x00000215839EA2B0> [label=2]
	<__main__.Node object at 0x0000021583A21470> [label=Survived]
	<__main__.Node object at 0x00000215839EA2B0> -> <__main__.Node object at 0x0000021583A21470> [label=0]
	<__main__.Node object at 0x0000021583A21588> [label=Survived]
	<__main__.Node object at 0x00000215839EA2B0> -> <__main__.Node object at 0x0000021583A21588> [label=3]
	<__main__.Node object at 0x0000021583A217F0> [label=Fare]
	<__main__.Node object at 0x00000215839EA2B0> -> <__main__.Node object at 0x0000021583A217F0> [label=1]
	<__main__.Node object at 0x0000021583A21780> [label=Embarked]
	<__main__.Node object at 0x0000021583A217F0> -> <__main__.Node object at 0x0000021583A21780> [label="upper class"]
	<__main__.Node object at 0x0000021583A21AC8> [label=Survived]
	<__main__.Node object at 0x0000021583A21780> -> <__main__.Node object at 0x0000021583A21AC8> [label=S]
	<__main__.Node object at 0x00000215839EAF28> [label=Survived]
	<__main__.Node object at 0x00000215839EA2B0> -> <__main__.Node object at 0x00000215839EAF28> [label=2]
	<__main__.Node object at 0x00000215839EA5C0> [label=Survived]
	<__main__.Node object at 0x00000215839F1668> -> <__main__.Node object at 0x00000215839EA5C0> [label=1]
	<__main__.Node object at 0x00000215839F1BA8> [label=Survived]
	<__main__.Node object at 0x00000215839F1A58> -> <__main__.Node object at 0x00000215839F1BA8> [label=teen]
	<__main__.Node object at 0x00000215839F18D0> [label=Death]
	<__main__.Node object at 0x00000215839F1A58> -> <__main__.Node object at 0x00000215839F18D0> [label=child]
	<__main__.Node object at 0x00000215829ACFD0> [label=Parch]
	<__main__.Node object at 0x00000215829AC5F8> -> <__main__.Node object at 0x00000215829ACFD0> [label=2]
	<__main__.Node object at 0x00000215839EAC50> [label=Survived]
	<__main__.Node object at 0x00000215829ACFD0> -> <__main__.Node object at 0x00000215839EAC50> [label=3]
	<__main__.Node object at 0x00000215839EAD68> [label=Survived]
	<__main__.Node object at 0x00000215829ACFD0> -> <__main__.Node object at 0x00000215839EAD68> [label=2]
	<__main__.Node object at 0x00000215839EA080> [label=Embarked]
	<__main__.Node object at 0x00000215829ACFD0> -> <__main__.Node object at 0x00000215839EA080> [label=0]
	<__main__.Node object at 0x0000021583A21358> [label=Age]
	<__main__.Node object at 0x00000215839EA080> -> <__main__.Node object at 0x0000021583A21358> [label=S]
	<__main__.Node object at 0x0000021583A21B38> [label=Survived]
	<__main__.Node object at 0x0000021583A21358> -> <__main__.Node object at 0x0000021583A21B38> [label=teen]
	<__main__.Node object at 0x0000021583A21CF8> [label=SibSp]
	<__main__.Node object at 0x0000021583A21358> -> <__main__.Node object at 0x0000021583A21CF8> [label=adults]
	<__main__.Node object at 0x0000021583A215C0> [label=Fare]
	<__main__.Node object at 0x0000021583A21CF8> -> <__main__.Node object at 0x0000021583A215C0> [label=0]
	<__main__.Node object at 0x00000215829641D0> [label=Survived]
	<__main__.Node object at 0x0000021583A215C0> -> <__main__.Node object at 0x00000215829641D0> [label="middle class"]
	<__main__.Node object at 0x0000021582964978> [label=Fare]
	<__main__.Node object at 0x0000021583A21CF8> -> <__main__.Node object at 0x0000021582964978> [label=1]
	<__main__.Node object at 0x0000021583A21F28> [label=Survived]
	<__main__.Node object at 0x0000021582964978> -> <__main__.Node object at 0x0000021583A21F28> [label="middle class"]
	<__main__.Node object at 0x0000021583A214A8> [label=Survived]
	<__main__.Node object at 0x00000215839EA080> -> <__main__.Node object at 0x0000021583A214A8> [label=C]
	<__main__.Node object at 0x0000021583A21B00> [label=Survived]
	<__main__.Node object at 0x00000215839EA080> -> <__main__.Node object at 0x0000021583A21B00> [label=Q]
	<__main__.Node object at 0x0000021583A211D0> [label=SibSp]
	<__main__.Node object at 0x00000215829ACFD0> -> <__main__.Node object at 0x0000021583A211D0> [label=1]
	<__main__.Node object at 0x0000021583A21550> [label=Age]
	<__main__.Node object at 0x0000021583A211D0> -> <__main__.Node object at 0x0000021583A21550> [label=1]
	<__main__.Node object at 0x0000021583A21D68> [label=Fare]
	<__main__.Node object at 0x0000021583A21550> -> <__main__.Node object at 0x0000021583A21D68> [label=adults]
	<__main__.Node object at 0x00000215839EA7B8> [label=Embarked]
	<__main__.Node object at 0x0000021583A21D68> -> <__main__.Node object at 0x00000215839EA7B8> [label="middle class"]
	<__main__.Node object at 0x00000215839EA908> [label=Survived]
	<__main__.Node object at 0x00000215839EA7B8> -> <__main__.Node object at 0x00000215839EA908> [label=S]
	<__main__.Node object at 0x0000021583A212B0> [label=Survived]
	<__main__.Node object at 0x0000021583A21550> -> <__main__.Node object at 0x0000021583A212B0> [label=child]
	<__main__.Node object at 0x0000021583A21CC0> [label=Survived]
	<__main__.Node object at 0x0000021583A211D0> -> <__main__.Node object at 0x0000021583A21CC0> [label=2]
	<__main__.Node object at 0x0000021583A219B0> [label=Survived]
	<__main__.Node object at 0x0000021583A211D0> -> <__main__.Node object at 0x0000021583A219B0> [label=0]
}
