digraph {
	<__main__.Node object at 0x00000168AAEFD5F8> [label=Sex]
	<__main__.Node object at 0x00000168B5CFA518> [label=Pclass]
	<__main__.Node object at 0x00000168AAEFD5F8> -> <__main__.Node object at 0x00000168B5CFA518> [label=male]
	<__main__.Node object at 0x00000168B5CFA940> [label=Age]
	<__main__.Node object at 0x00000168B5CFA518> -> <__main__.Node object at 0x00000168B5CFA940> [label=2]
	<__main__.Node object at 0x00000168B5CFA550> [label=Parch]
	<__main__.Node object at 0x00000168B5CFA940> -> <__main__.Node object at 0x00000168B5CFA550> [label=adults]
	<__main__.Node object at 0x00000168B5CDB048> [label=Fare]
	<__main__.Node object at 0x00000168B5CFA550> -> <__main__.Node object at 0x00000168B5CDB048> [label=0]
	<__main__.Node object at 0x00000168B5CFAD30> [label=Embarked]
	<__main__.Node object at 0x00000168B5CDB048> -> <__main__.Node object at 0x00000168B5CFAD30> [label="middle class"]
	<__main__.Node object at 0x00000168B5CDB978> [label=SibSp]
	<__main__.Node object at 0x00000168B5CFAD30> -> <__main__.Node object at 0x00000168B5CDB978> [label=S]
	<__main__.Node object at 0x00000168B5CDB160> [label=Death]
	<__main__.Node object at 0x00000168B5CDB978> -> <__main__.Node object at 0x00000168B5CDB160> [label=1]
	<__main__.Node object at 0x00000168B5CDB550> [label=Death]
	<__main__.Node object at 0x00000168B5CDB978> -> <__main__.Node object at 0x00000168B5CDB550> [label=0]
	<__main__.Node object at 0x00000168B5CDB208> [label=SibSp]
	<__main__.Node object at 0x00000168B5CFAD30> -> <__main__.Node object at 0x00000168B5CDB208> [label=C]
	<__main__.Node object at 0x00000168B5CDB0B8> [label=Death]
	<__main__.Node object at 0x00000168B5CDB208> -> <__main__.Node object at 0x00000168B5CDB0B8> [label=0]
	<__main__.Node object at 0x00000168B5CDB358> [label=Death]
	<__main__.Node object at 0x00000168B5CDB208> -> <__main__.Node object at 0x00000168B5CDB358> [label=1]
	<__main__.Node object at 0x00000168B4C75F60> [label=Death]
	<__main__.Node object at 0x00000168B5CDB048> -> <__main__.Node object at 0x00000168B4C75F60> [label=poor]
	<__main__.Node object at 0x00000168B5C91F98> [label=Death]
	<__main__.Node object at 0x00000168B5CDB048> -> <__main__.Node object at 0x00000168B5C91F98> [label="upper class"]
	<__main__.Node object at 0x00000168B5CFA860> [label=Death]
	<__main__.Node object at 0x00000168B5CFA550> -> <__main__.Node object at 0x00000168B5CFA860> [label=2]
	<__main__.Node object at 0x00000168B5C91DD8> [label=Death]
	<__main__.Node object at 0x00000168B5CFA550> -> <__main__.Node object at 0x00000168B5C91DD8> [label=1]
	<__main__.Node object at 0x00000168B4723320> [label=Death]
	<__main__.Node object at 0x00000168B5CFA940> -> <__main__.Node object at 0x00000168B4723320> [label=teen]
	<__main__.Node object at 0x00000168B5C91BA8> [label=Survived]
	<__main__.Node object at 0x00000168B5CFA940> -> <__main__.Node object at 0x00000168B5C91BA8> [label=child]
	<__main__.Node object at 0x00000168B5CFAF98> [label=Death]
	<__main__.Node object at 0x00000168B5CFA940> -> <__main__.Node object at 0x00000168B5CFAF98> [label=elderly]
	<__main__.Node object at 0x00000168B5CFAC50> [label=SibSp]
	<__main__.Node object at 0x00000168B5CFA518> -> <__main__.Node object at 0x00000168B5CFAC50> [label=3]
	<__main__.Node object at 0x00000168B5CFAEB8> [label=Death]
	<__main__.Node object at 0x00000168B5CFAC50> -> <__main__.Node object at 0x00000168B5CFAEB8> [label=8]
	<__main__.Node object at 0x00000168B5CFAEF0> [label=Fare]
	<__main__.Node object at 0x00000168B5CFAC50> -> <__main__.Node object at 0x00000168B5CFAEF0> [label=0]
	<__main__.Node object at 0x00000168B5CFAF60> [label=Age]
	<__main__.Node object at 0x00000168B5CFAEF0> -> <__main__.Node object at 0x00000168B5CFAF60> [label=poor]
	<__main__.Node object at 0x00000168B5CDB390> [label=Parch]
	<__main__.Node object at 0x00000168B5CFAF60> -> <__main__.Node object at 0x00000168B5CDB390> [label=adults]
	<__main__.Node object at 0x00000168B5CDBBA8> [label=Embarked]
	<__main__.Node object at 0x00000168B5CDB390> -> <__main__.Node object at 0x00000168B5CDBBA8> [label=0]
	<__main__.Node object at 0x00000168B5CDBCF8> [label=Death]
	<__main__.Node object at 0x00000168B5CDBBA8> -> <__main__.Node object at 0x00000168B5CDBCF8> [label=C]
	<__main__.Node object at 0x00000168B5CDBC88> [label=Death]
	<__main__.Node object at 0x00000168B5CDBBA8> -> <__main__.Node object at 0x00000168B5CDBC88> [label=S]
	<__main__.Node object at 0x00000168B5CDBD68> [label=Death]
	<__main__.Node object at 0x00000168B5CDBBA8> -> <__main__.Node object at 0x00000168B5CDBD68> [label=Q]
	<__main__.Node object at 0x00000168B5CDB898> [label=Death]
	<__main__.Node object at 0x00000168B5CDB390> -> <__main__.Node object at 0x00000168B5CDB898> [label=1]
	<__main__.Node object at 0x00000168B5CDBA20> [label=Parch]
	<__main__.Node object at 0x00000168B5CFAF60> -> <__main__.Node object at 0x00000168B5CDBA20> [label=teen]
	<__main__.Node object at 0x00000168B5CDB630> [label=Embarked]
	<__main__.Node object at 0x00000168B5CDBA20> -> <__main__.Node object at 0x00000168B5CDB630> [label=0]
	<__main__.Node object at 0x00000168B5CDBE10> [label=Death]
	<__main__.Node object at 0x00000168B5CDB630> -> <__main__.Node object at 0x00000168B5CDBE10> [label=S]
	<__main__.Node object at 0x00000168B5CDBC50> [label=Death]
	<__main__.Node object at 0x00000168B5CFAF60> -> <__main__.Node object at 0x00000168B5CDBC50> [label=elderly]
	<__main__.Node object at 0x00000168B5CDB2B0> [label=Age]
	<__main__.Node object at 0x00000168B5CFAEF0> -> <__main__.Node object at 0x00000168B5CDB2B0> [label="middle class"]
	<__main__.Node object at 0x00000168B5CDB908> [label=Death]
	<__main__.Node object at 0x00000168B5CDB2B0> -> <__main__.Node object at 0x00000168B5CDB908> [label=adults]
	<__main__.Node object at 0x00000168B5CDB828> [label=Parch]
	<__main__.Node object at 0x00000168B5CDB2B0> -> <__main__.Node object at 0x00000168B5CDB828> [label=child]
	<__main__.Node object at 0x00000168B5CDB128> [label=Death]
	<__main__.Node object at 0x00000168B5CDB828> -> <__main__.Node object at 0x00000168B5CDB128> [label=0]
	<__main__.Node object at 0x00000168B5CDBB38> [label=Survived]
	<__main__.Node object at 0x00000168B5CDB828> -> <__main__.Node object at 0x00000168B5CDBB38> [label=1]
	<__main__.Node object at 0x00000168B5CDB1D0> [label=Age]
	<__main__.Node object at 0x00000168B5CFAEF0> -> <__main__.Node object at 0x00000168B5CDB1D0> [label="upper class"]
	<__main__.Node object at 0x00000168B5CDB470> [label=Parch]
	<__main__.Node object at 0x00000168B5CDB1D0> -> <__main__.Node object at 0x00000168B5CDB470> [label=adults]
	<__main__.Node object at 0x00000168B5CDBDA0> [label=Embarked]
	<__main__.Node object at 0x00000168B5CDB470> -> <__main__.Node object at 0x00000168B5CDBDA0> [label=0]
	<__main__.Node object at 0x00000168B5CADF28> [label=Survived]
	<__main__.Node object at 0x00000168B5CDBDA0> -> <__main__.Node object at 0x00000168B5CADF28> [label=S]
	<__main__.Node object at 0x00000168B5C91FD0> [label=Age]
	<__main__.Node object at 0x00000168B5CFAC50> -> <__main__.Node object at 0x00000168B5C91FD0> [label=1]
	<__main__.Node object at 0x00000168B5CDBB00> [label=Embarked]
	<__main__.Node object at 0x00000168B5C91FD0> -> <__main__.Node object at 0x00000168B5CDBB00> [label=adults]
	<__main__.Node object at 0x00000168B5CDB5C0> [label=Fare]
	<__main__.Node object at 0x00000168B5CDBB00> -> <__main__.Node object at 0x00000168B5CDB5C0> [label=S]
	<__main__.Node object at 0x00000168B5CADCC0> [label=Death]
	<__main__.Node object at 0x00000168B5CDB5C0> -> <__main__.Node object at 0x00000168B5CADCC0> [label="middle class"]
	<__main__.Node object at 0x00000168B5CADA90> [label=Parch]
	<__main__.Node object at 0x00000168B5CDB5C0> -> <__main__.Node object at 0x00000168B5CADA90> [label=poor]
	<__main__.Node object at 0x00000168B5CADE48> [label=Death]
	<__main__.Node object at 0x00000168B5CADA90> -> <__main__.Node object at 0x00000168B5CADE48> [label=0]
	<__main__.Node object at 0x00000168B5CDBFD0> [label=Parch]
	<__main__.Node object at 0x00000168B5CDBB00> -> <__main__.Node object at 0x00000168B5CDBFD0> [label=C]
	<__main__.Node object at 0x00000168B5CDB2E8> [label=Survived]
	<__main__.Node object at 0x00000168B5CDBFD0> -> <__main__.Node object at 0x00000168B5CDB2E8> [label=1]
	<__main__.Node object at 0x00000168B5CDBC18> [label=Death]
	<__main__.Node object at 0x00000168B5CDBFD0> -> <__main__.Node object at 0x00000168B5CDBC18> [label=0]
	<__main__.Node object at 0x00000168B5CDB3C8> [label=Death]
	<__main__.Node object at 0x00000168B5CDBB00> -> <__main__.Node object at 0x00000168B5CDB3C8> [label=Q]
	<__main__.Node object at 0x00000168B5CDB748> [label=Death]
	<__main__.Node object at 0x00000168B5C91FD0> -> <__main__.Node object at 0x00000168B5CDB748> [label=teen]
	<__main__.Node object at 0x00000168B5CDB780> [label=Survived]
	<__main__.Node object at 0x00000168B5C91FD0> -> <__main__.Node object at 0x00000168B5CDB780> [label=child]
	<__main__.Node object at 0x00000168B5CFA470> [label=Death]
	<__main__.Node object at 0x00000168B5CFAC50> -> <__main__.Node object at 0x00000168B5CFA470> [label=3]
	<__main__.Node object at 0x00000168B5CFA358> [label=Embarked]
	<__main__.Node object at 0x00000168B5CFAC50> -> <__main__.Node object at 0x00000168B5CFA358> [label=2]
	<__main__.Node object at 0x00000168B5CDBD30> [label=Death]
	<__main__.Node object at 0x00000168B5CFA358> -> <__main__.Node object at 0x00000168B5CDBD30> [label=S]
	<__main__.Node object at 0x00000168B5CDB940> [label=Survived]
	<__main__.Node object at 0x00000168B5CFA358> -> <__main__.Node object at 0x00000168B5CDB940> [label=Q]
	<__main__.Node object at 0x00000168B5C91F60> [label=Death]
	<__main__.Node object at 0x00000168B5CFAC50> -> <__main__.Node object at 0x00000168B5C91F60> [label=5]
	<__main__.Node object at 0x00000168B5C91F28> [label=Parch]
	<__main__.Node object at 0x00000168B5CFAC50> -> <__main__.Node object at 0x00000168B5C91F28> [label=4]
	<__main__.Node object at 0x00000168B5CDB518> [label=Age]
	<__main__.Node object at 0x00000168B5C91F28> -> <__main__.Node object at 0x00000168B5CDB518> [label=2]
	<__main__.Node object at 0x00000168B5CADB00> [label=Fare]
	<__main__.Node object at 0x00000168B5CDB518> -> <__main__.Node object at 0x00000168B5CADB00> [label=child]
	<__main__.Node object at 0x00000168B5CAD5C0> [label=Embarked]
	<__main__.Node object at 0x00000168B5CADB00> -> <__main__.Node object at 0x00000168B5CAD5C0> [label="middle class"]
	<__main__.Node object at 0x00000168B5CAD2E8> [label=Death]
	<__main__.Node object at 0x00000168B5CAD5C0> -> <__main__.Node object at 0x00000168B5CAD2E8> [label=S]
	<__main__.Node object at 0x00000168B5CDB710> [label=Death]
	<__main__.Node object at 0x00000168B5C91F28> -> <__main__.Node object at 0x00000168B5CDB710> [label=1]
	<__main__.Node object at 0x00000168B5CFA8D0> [label=Age]
	<__main__.Node object at 0x00000168B5CFA518> -> <__main__.Node object at 0x00000168B5CFA8D0> [label=1]
	<__main__.Node object at 0x00000168B5CDBE80> [label=SibSp]
	<__main__.Node object at 0x00000168B5CFA8D0> -> <__main__.Node object at 0x00000168B5CDBE80> [label=adults]
	<__main__.Node object at 0x00000168B5CADF60> [label=Fare]
	<__main__.Node object at 0x00000168B5CDBE80> -> <__main__.Node object at 0x00000168B5CADF60> [label=0]
	<__main__.Node object at 0x00000168B5CAD940> [label=Embarked]
	<__main__.Node object at 0x00000168B5CADF60> -> <__main__.Node object at 0x00000168B5CAD940> [label="middle class"]
	<__main__.Node object at 0x00000168B5CAD240> [label=Parch]
	<__main__.Node object at 0x00000168B5CAD940> -> <__main__.Node object at 0x00000168B5CAD240> [label=C]
	<__main__.Node object at 0x00000168B5CADCF8> [label=Death]
	<__main__.Node object at 0x00000168B5CAD240> -> <__main__.Node object at 0x00000168B5CADCF8> [label=0]
	<__main__.Node object at 0x00000168B5CAD080> [label=Parch]
	<__main__.Node object at 0x00000168B5CAD940> -> <__main__.Node object at 0x00000168B5CAD080> [label=S]
	<__main__.Node object at 0x00000168B5CAD358> [label=Death]
	<__main__.Node object at 0x00000168B5CAD080> -> <__main__.Node object at 0x00000168B5CAD358> [label=0]
	<__main__.Node object at 0x00000168B5CADE80> [label=Death]
	<__main__.Node object at 0x00000168B5CADF60> -> <__main__.Node object at 0x00000168B5CADE80> [label=poor]
	<__main__.Node object at 0x00000168B5CAD2B0> [label=Embarked]
	<__main__.Node object at 0x00000168B5CADF60> -> <__main__.Node object at 0x00000168B5CAD2B0> [label="upper class"]
	<__main__.Node object at 0x00000168B5CAD400> [label=Death]
	<__main__.Node object at 0x00000168B5CAD2B0> -> <__main__.Node object at 0x00000168B5CAD400> [label=S]
	<__main__.Node object at 0x00000168B5CAD438> [label=Parch]
	<__main__.Node object at 0x00000168B5CAD2B0> -> <__main__.Node object at 0x00000168B5CAD438> [label=C]
	<__main__.Node object at 0x00000168B5CAD128> [label=Death]
	<__main__.Node object at 0x00000168B5CAD438> -> <__main__.Node object at 0x00000168B5CAD128> [label=0]
	<__main__.Node object at 0x00000168B5CAD390> [label=Survived]
	<__main__.Node object at 0x00000168B5CAD438> -> <__main__.Node object at 0x00000168B5CAD390> [label=1]
	<__main__.Node object at 0x00000168B5CADFD0> [label=Death]
	<__main__.Node object at 0x00000168B5CAD438> -> <__main__.Node object at 0x00000168B5CADFD0> [label=2]
	<__main__.Node object at 0x00000168B5CADDA0> [label=Death]
	<__main__.Node object at 0x00000168B5CDBE80> -> <__main__.Node object at 0x00000168B5CADDA0> [label=2]
	<__main__.Node object at 0x00000168B5CADC88> [label=Parch]
	<__main__.Node object at 0x00000168B5CDBE80> -> <__main__.Node object at 0x00000168B5CADC88> [label=1]
	<__main__.Node object at 0x00000168B5CADD30> [label=Embarked]
	<__main__.Node object at 0x00000168B5CADC88> -> <__main__.Node object at 0x00000168B5CADD30> [label=0]
	<__main__.Node object at 0x00000168B5CAD7B8> [label=Fare]
	<__main__.Node object at 0x00000168B5CADD30> -> <__main__.Node object at 0x00000168B5CAD7B8> [label=C]
	<__main__.Node object at 0x00000168B5CDB080> [label=Survived]
	<__main__.Node object at 0x00000168B5CAD7B8> -> <__main__.Node object at 0x00000168B5CDB080> [label="upper class"]
	<__main__.Node object at 0x00000168B5CAD748> [label=Fare]
	<__main__.Node object at 0x00000168B5CADD30> -> <__main__.Node object at 0x00000168B5CAD748> [label=S]
	<__main__.Node object at 0x00000168B5CAD588> [label=Death]
	<__main__.Node object at 0x00000168B5CAD748> -> <__main__.Node object at 0x00000168B5CAD588> [label="upper class"]
	<__main__.Node object at 0x00000168B5CAD6A0> [label=Survived]
	<__main__.Node object at 0x00000168B5CADC88> -> <__main__.Node object at 0x00000168B5CAD6A0> [label=2]
	<__main__.Node object at 0x00000168B5CAD278> [label=Embarked]
	<__main__.Node object at 0x00000168B5CADC88> -> <__main__.Node object at 0x00000168B5CAD278> [label=1]
	<__main__.Node object at 0x00000168B5CADC50> [label=Fare]
	<__main__.Node object at 0x00000168B5CAD278> -> <__main__.Node object at 0x00000168B5CADC50> [label=C]
	<__main__.Node object at 0x00000168B5CDBA90> [label=Survived]
	<__main__.Node object at 0x00000168B5CADC50> -> <__main__.Node object at 0x00000168B5CDBA90> [label="upper class"]
	<__main__.Node object at 0x00000168B5CAD9E8> [label=Survived]
	<__main__.Node object at 0x00000168B5CAD278> -> <__main__.Node object at 0x00000168B5CAD9E8> [label=S]
	<__main__.Node object at 0x00000168B5CAD160> [label=Death]
	<__main__.Node object at 0x00000168B5CADC88> -> <__main__.Node object at 0x00000168B5CAD160> [label=4]
	<__main__.Node object at 0x00000168B5C91198> [label=Death]
	<__main__.Node object at 0x00000168B5CDBE80> -> <__main__.Node object at 0x00000168B5C91198> [label=3]
	<__main__.Node object at 0x00000168B5CAD978> [label=Survived]
	<__main__.Node object at 0x00000168B5CFA8D0> -> <__main__.Node object at 0x00000168B5CAD978> [label=child]
	<__main__.Node object at 0x00000168B5CAD7F0> [label=Death]
	<__main__.Node object at 0x00000168B5CFA8D0> -> <__main__.Node object at 0x00000168B5CAD7F0> [label=elderly]
	<__main__.Node object at 0x00000168B5CAD908> [label=SibSp]
	<__main__.Node object at 0x00000168B5CFA8D0> -> <__main__.Node object at 0x00000168B5CAD908> [label=teen]
	<__main__.Node object at 0x00000168B5CAD710> [label=Death]
	<__main__.Node object at 0x00000168B5CAD908> -> <__main__.Node object at 0x00000168B5CAD710> [label=1]
	<__main__.Node object at 0x00000168B5CADEB8> [label=Survived]
	<__main__.Node object at 0x00000168B5CAD908> -> <__main__.Node object at 0x00000168B5CADEB8> [label=0]
	<__main__.Node object at 0x00000168B5C91780> [label=Pclass]
	<__main__.Node object at 0x00000168AAEFD5F8> -> <__main__.Node object at 0x00000168B5C91780> [label=female]
	<__main__.Node object at 0x00000168B5CAD048> [label=SibSp]
	<__main__.Node object at 0x00000168B5C91780> -> <__main__.Node object at 0x00000168B5CAD048> [label=3]
	<__main__.Node object at 0x00000168B5CDBAC8> [label=Parch]
	<__main__.Node object at 0x00000168B5CAD048> -> <__main__.Node object at 0x00000168B5CDBAC8> [label=1]
	<__main__.Node object at 0x00000168B5CFABA8> [label=Embarked]
	<__main__.Node object at 0x00000168B5CDBAC8> -> <__main__.Node object at 0x00000168B5CFABA8> [label=0]
	<__main__.Node object at 0x00000168B5CFA4E0> [label=Fare]
	<__main__.Node object at 0x00000168B5CFABA8> -> <__main__.Node object at 0x00000168B5CFA4E0> [label=S]
	<__main__.Node object at 0x00000168B4C93A20> [label=Age]
	<__main__.Node object at 0x00000168B5CFA4E0> -> <__main__.Node object at 0x00000168B4C93A20> [label=poor]
	<__main__.Node object at 0x00000168B4C93BE0> [label=Death]
	<__main__.Node object at 0x00000168B4C93A20> -> <__main__.Node object at 0x00000168B4C93BE0> [label=adults]
	<__main__.Node object at 0x00000168B4C93CC0> [label=Age]
	<__main__.Node object at 0x00000168B5CFA4E0> -> <__main__.Node object at 0x00000168B4C93CC0> [label="middle class"]
	<__main__.Node object at 0x00000168B4C93B38> [label=Death]
	<__main__.Node object at 0x00000168B4C93CC0> -> <__main__.Node object at 0x00000168B4C93B38> [label=adults]
	<__main__.Node object at 0x00000168B5CFAE48> [label=Survived]
	<__main__.Node object at 0x00000168B5CFABA8> -> <__main__.Node object at 0x00000168B5CFAE48> [label=Q]
	<__main__.Node object at 0x00000168B5CFA5F8> [label=Age]
	<__main__.Node object at 0x00000168B5CFABA8> -> <__main__.Node object at 0x00000168B5CFA5F8> [label=C]
	<__main__.Node object at 0x00000168B4C93128> [label=Fare]
	<__main__.Node object at 0x00000168B5CFA5F8> -> <__main__.Node object at 0x00000168B4C93128> [label=teen]
	<__main__.Node object at 0x00000168B4C932B0> [label=Survived]
	<__main__.Node object at 0x00000168B4C93128> -> <__main__.Node object at 0x00000168B4C932B0> [label="middle class"]
	<__main__.Node object at 0x00000168B5CFA9E8> [label=Embarked]
	<__main__.Node object at 0x00000168B5CDBAC8> -> <__main__.Node object at 0x00000168B5CFA9E8> [label=1]
	<__main__.Node object at 0x00000168B5CFA978> [label=Age]
	<__main__.Node object at 0x00000168B5CFA9E8> -> <__main__.Node object at 0x00000168B5CFA978> [label=S]
	<__main__.Node object at 0x00000168B4C93B70> [label=Fare]
	<__main__.Node object at 0x00000168B5CFA978> -> <__main__.Node object at 0x00000168B4C93B70> [label=adults]
	<__main__.Node object at 0x00000168B4C93160> [label=Death]
	<__main__.Node object at 0x00000168B4C93B70> -> <__main__.Node object at 0x00000168B4C93160> [label="middle class"]
	<__main__.Node object at 0x00000168B4C93A58> [label=Survived]
	<__main__.Node object at 0x00000168B5CFA978> -> <__main__.Node object at 0x00000168B4C93A58> [label=child]
	<__main__.Node object at 0x00000168B5CFAB70> [label=Death]
	<__main__.Node object at 0x00000168B5CFA9E8> -> <__main__.Node object at 0x00000168B5CFAB70> [label=Q]
	<__main__.Node object at 0x00000168B5CFAA58> [label=Age]
	<__main__.Node object at 0x00000168B5CFA9E8> -> <__main__.Node object at 0x00000168B5CFAA58> [label=C]
	<__main__.Node object at 0x00000168AD344358> [label=Survived]
	<__main__.Node object at 0x00000168B5CFAA58> -> <__main__.Node object at 0x00000168AD344358> [label=adults]
	<__main__.Node object at 0x00000168B4C93B00> [label=Death]
	<__main__.Node object at 0x00000168B5CFAA58> -> <__main__.Node object at 0x00000168B4C93B00> [label=child]
	<__main__.Node object at 0x00000168B5CFACC0> [label=Death]
	<__main__.Node object at 0x00000168B5CDBAC8> -> <__main__.Node object at 0x00000168B5CFACC0> [label=6]
	<__main__.Node object at 0x00000168B45D2D68> [label=Survived]
	<__main__.Node object at 0x00000168B5CDBAC8> -> <__main__.Node object at 0x00000168B45D2D68> [label=5]
	<__main__.Node object at 0x00000168B5CFAF28> [label=Death]
	<__main__.Node object at 0x00000168B5CDBAC8> -> <__main__.Node object at 0x00000168B5CFAF28> [label=3]
	<__main__.Node object at 0x00000168B5CFACF8> [label=Death]
	<__main__.Node object at 0x00000168B5CDBAC8> -> <__main__.Node object at 0x00000168B5CFACF8> [label=2]
	<__main__.Node object at 0x00000168B5CFADA0> [label=Death]
	<__main__.Node object at 0x00000168B5CDBAC8> -> <__main__.Node object at 0x00000168B5CFADA0> [label=4]
	<__main__.Node object at 0x00000168B5CFA898> [label=Age]
	<__main__.Node object at 0x00000168B5CAD048> -> <__main__.Node object at 0x00000168B5CFA898> [label=4]
	<__main__.Node object at 0x00000168B5CDB5F8> [label=Parch]
	<__main__.Node object at 0x00000168B5CFA898> -> <__main__.Node object at 0x00000168B5CDB5F8> [label=child]
	<__main__.Node object at 0x00000168B5CDB668> [label=Fare]
	<__main__.Node object at 0x00000168B5CDB5F8> -> <__main__.Node object at 0x00000168B5CDB668> [label=2]
	<__main__.Node object at 0x00000168B5CAFE48> [label=Embarked]
	<__main__.Node object at 0x00000168B5CDB668> -> <__main__.Node object at 0x00000168B5CAFE48> [label="middle class"]
	<__main__.Node object at 0x00000168B4C939B0> [label=Death]
	<__main__.Node object at 0x00000168B5CAFE48> -> <__main__.Node object at 0x00000168B4C939B0> [label=S]
	<__main__.Node object at 0x00000168B4C93208> [label=Survived]
	<__main__.Node object at 0x00000168B5CFA898> -> <__main__.Node object at 0x00000168B4C93208> [label=teen]
	<__main__.Node object at 0x00000168B4C934A8> [label=Parch]
	<__main__.Node object at 0x00000168B5CAD048> -> <__main__.Node object at 0x00000168B4C934A8> [label=0]
	<__main__.Node object at 0x00000168B4C938D0> [label=Embarked]
	<__main__.Node object at 0x00000168B4C934A8> -> <__main__.Node object at 0x00000168B4C938D0> [label=2]
	<__main__.Node object at 0x00000168B4C93BA8> [label=Survived]
	<__main__.Node object at 0x00000168B4C938D0> -> <__main__.Node object at 0x00000168B4C93BA8> [label=S]
	<__main__.Node object at 0x00000168B5CFA6D8> [label=Age]
	<__main__.Node object at 0x00000168B4C938D0> -> <__main__.Node object at 0x00000168B5CFA6D8> [label=C]
	<__main__.Node object at 0x00000168B5CFA710> [label=Survived]
	<__main__.Node object at 0x00000168B5CFA6D8> -> <__main__.Node object at 0x00000168B5CFA710> [label=child]
	<__main__.Node object at 0x00000168B5CFAC88> [label=Fare]
	<__main__.Node object at 0x00000168B5CFA6D8> -> <__main__.Node object at 0x00000168B5CFAC88> [label=adults]
	<__main__.Node object at 0x00000168B5CDB4A8> [label=Survived]
	<__main__.Node object at 0x00000168B5CFAC88> -> <__main__.Node object at 0x00000168B5CDB4A8> [label="middle class"]
	<__main__.Node object at 0x00000168B5CFADD8> [label=Death]
	<__main__.Node object at 0x00000168B4C938D0> -> <__main__.Node object at 0x00000168B5CFADD8> [label=Q]
	<__main__.Node object at 0x00000168B4C93DD8> [label=Embarked]
	<__main__.Node object at 0x00000168B4C934A8> -> <__main__.Node object at 0x00000168B4C93DD8> [label=0]
	<__main__.Node object at 0x00000168B4C93EB8> [label=Age]
	<__main__.Node object at 0x00000168B4C93DD8> -> <__main__.Node object at 0x00000168B4C93EB8> [label=S]
	<__main__.Node object at 0x00000168B5CAD828> [label=Fare]
	<__main__.Node object at 0x00000168B4C93EB8> -> <__main__.Node object at 0x00000168B5CAD828> [label=adults]
	<__main__.Node object at 0x00000168B5CAFC18> [label=Death]
	<__main__.Node object at 0x00000168B5CAD828> -> <__main__.Node object at 0x00000168B5CAFC18> [label=poor]
	<__main__.Node object at 0x00000168B5CAFE80> [label=Survived]
	<__main__.Node object at 0x00000168B5CAD828> -> <__main__.Node object at 0x00000168B5CAFE80> [label="middle class"]
	<__main__.Node object at 0x00000168B5CADD68> [label=Survived]
	<__main__.Node object at 0x00000168B4C93EB8> -> <__main__.Node object at 0x00000168B5CADD68> [label=child]
	<__main__.Node object at 0x00000168B4C932E8> [label=Age]
	<__main__.Node object at 0x00000168B4C93DD8> -> <__main__.Node object at 0x00000168B4C932E8> [label=Q]
	<__main__.Node object at 0x00000168B5CAD860> [label=Fare]
	<__main__.Node object at 0x00000168B4C932E8> -> <__main__.Node object at 0x00000168B5CAD860> [label=adults]
	<__main__.Node object at 0x00000168B5CAFEF0> [label=Survived]
	<__main__.Node object at 0x00000168B5CAD860> -> <__main__.Node object at 0x00000168B5CAFEF0> [label=poor]
	<__main__.Node object at 0x00000168B5CFA9B0> [label=Survived]
	<__main__.Node object at 0x00000168B4C932E8> -> <__main__.Node object at 0x00000168B5CFA9B0> [label=teen]
	<__main__.Node object at 0x00000168B5CADE10> [label=Fare]
	<__main__.Node object at 0x00000168B4C93DD8> -> <__main__.Node object at 0x00000168B5CADE10> [label=C]
	<__main__.Node object at 0x00000168B5CDB0F0> [label=Survived]
	<__main__.Node object at 0x00000168B5CADE10> -> <__main__.Node object at 0x00000168B5CDB0F0> [label=poor]
	<__main__.Node object at 0x00000168B5CDBDD8> [label=Death]
	<__main__.Node object at 0x00000168B5CADE10> -> <__main__.Node object at 0x00000168B5CDBDD8> [label="middle class"]
	<__main__.Node object at 0x00000168B5CFAAC8> [label=Embarked]
	<__main__.Node object at 0x00000168B4C934A8> -> <__main__.Node object at 0x00000168B5CFAAC8> [label=1]
	<__main__.Node object at 0x00000168B4C93390> [label=Death]
	<__main__.Node object at 0x00000168B5CFAAC8> -> <__main__.Node object at 0x00000168B4C93390> [label=C]
	<__main__.Node object at 0x00000168B4C939E8> [label=Age]
	<__main__.Node object at 0x00000168B5CFAAC8> -> <__main__.Node object at 0x00000168B4C939E8> [label=S]
	<__main__.Node object at 0x00000168B5CAF198> [label=Fare]
	<__main__.Node object at 0x00000168B4C939E8> -> <__main__.Node object at 0x00000168B5CAF198> [label=child]
	<__main__.Node object at 0x00000168B5D23240> [label=Survived]
	<__main__.Node object at 0x00000168B5CAF198> -> <__main__.Node object at 0x00000168B5D23240> [label="middle class"]
	<__main__.Node object at 0x00000168B5CAF940> [label=Survived]
	<__main__.Node object at 0x00000168B4C939E8> -> <__main__.Node object at 0x00000168B5CAF940> [label=adults]
	<__main__.Node object at 0x00000168B5CAF1D0> [label=Survived]
	<__main__.Node object at 0x00000168B4C939E8> -> <__main__.Node object at 0x00000168B5CAF1D0> [label=teen]
	<__main__.Node object at 0x00000168B5CDB8D0> [label=Death]
	<__main__.Node object at 0x00000168B4C934A8> -> <__main__.Node object at 0x00000168B5CDB8D0> [label=4]
	<__main__.Node object at 0x00000168B5CDB588> [label=Death]
	<__main__.Node object at 0x00000168B4C934A8> -> <__main__.Node object at 0x00000168B5CDB588> [label=5]
	<__main__.Node object at 0x00000168B5CFA780> [label=Parch]
	<__main__.Node object at 0x00000168B5CAD048> -> <__main__.Node object at 0x00000168B5CFA780> [label=3]
	<__main__.Node object at 0x00000168B4C93748> [label=Survived]
	<__main__.Node object at 0x00000168B5CFA780> -> <__main__.Node object at 0x00000168B4C93748> [label=0]
	<__main__.Node object at 0x00000168B4C937B8> [label=Death]
	<__main__.Node object at 0x00000168B5CFA780> -> <__main__.Node object at 0x00000168B4C937B8> [label=1]
	<__main__.Node object at 0x00000168B4C93CF8> [label=Death]
	<__main__.Node object at 0x00000168B5CFA780> -> <__main__.Node object at 0x00000168B4C93CF8> [label=2]
	<__main__.Node object at 0x00000168B5CFAE80> [label=Embarked]
	<__main__.Node object at 0x00000168B5CAD048> -> <__main__.Node object at 0x00000168B5CFAE80> [label=2]
	<__main__.Node object at 0x00000168B4C93C88> [label=Death]
	<__main__.Node object at 0x00000168B5CFAE80> -> <__main__.Node object at 0x00000168B4C93C88> [label=S]
	<__main__.Node object at 0x00000168B4C93320> [label=Survived]
	<__main__.Node object at 0x00000168B5CFAE80> -> <__main__.Node object at 0x00000168B4C93320> [label=C]
	<__main__.Node object at 0x00000168B4C934E0> [label=Survived]
	<__main__.Node object at 0x00000168B5CFAE80> -> <__main__.Node object at 0x00000168B4C934E0> [label=Q]
	<__main__.Node object at 0x00000168B5CADBE0> [label=Death]
	<__main__.Node object at 0x00000168B5CAD048> -> <__main__.Node object at 0x00000168B5CADBE0> [label=8]
	<__main__.Node object at 0x00000168B5CAD198> [label=Death]
	<__main__.Node object at 0x00000168B5CAD048> -> <__main__.Node object at 0x00000168B5CAD198> [label=5]
	<__main__.Node object at 0x00000168B5CAD320> [label=Age]
	<__main__.Node object at 0x00000168B5C91780> -> <__main__.Node object at 0x00000168B5CAD320> [label=1]
	<__main__.Node object at 0x00000168B5CDB4E0> [label=Parch]
	<__main__.Node object at 0x00000168B5CAD320> -> <__main__.Node object at 0x00000168B5CDB4E0> [label=adults]
	<__main__.Node object at 0x00000168B5CAF208> [label=Fare]
	<__main__.Node object at 0x00000168B5CDB4E0> -> <__main__.Node object at 0x00000168B5CAF208> [label=0]
	<__main__.Node object at 0x00000168B5D235C0> [label=Survived]
	<__main__.Node object at 0x00000168B5CAF208> -> <__main__.Node object at 0x00000168B5D235C0> [label="upper class"]
	<__main__.Node object at 0x00000168B5D231D0> [label=Embarked]
	<__main__.Node object at 0x00000168B5CAF208> -> <__main__.Node object at 0x00000168B5D231D0> [label="middle class"]
	<__main__.Node object at 0x00000168B5D236D8> [label=SibSp]
	<__main__.Node object at 0x00000168B5D231D0> -> <__main__.Node object at 0x00000168B5D236D8> [label=C]
	<__main__.Node object at 0x00000168B5D238D0> [label=Survived]
	<__main__.Node object at 0x00000168B5D236D8> -> <__main__.Node object at 0x00000168B5D238D0> [label=0]
	<__main__.Node object at 0x00000168B5D239E8> [label=Survived]
	<__main__.Node object at 0x00000168B5D236D8> -> <__main__.Node object at 0x00000168B5D239E8> [label=1]
	<__main__.Node object at 0x00000168B5D23470> [label=Survived]
	<__main__.Node object at 0x00000168B5D231D0> -> <__main__.Node object at 0x00000168B5D23470> [label=S]
	<__main__.Node object at 0x00000168B5CAFA90> [label=Survived]
	<__main__.Node object at 0x00000168B5CDB4E0> -> <__main__.Node object at 0x00000168B5CAFA90> [label=1]
	<__main__.Node object at 0x00000168B5CAF0F0> [label=SibSp]
	<__main__.Node object at 0x00000168B5CDB4E0> -> <__main__.Node object at 0x00000168B5CAF0F0> [label=2]
	<__main__.Node object at 0x00000168B5D23198> [label=Survived]
	<__main__.Node object at 0x00000168B5CAF0F0> -> <__main__.Node object at 0x00000168B5D23198> [label=0]
	<__main__.Node object at 0x00000168B5D23668> [label=Survived]
	<__main__.Node object at 0x00000168B5CAF0F0> -> <__main__.Node object at 0x00000168B5D23668> [label=2]
	<__main__.Node object at 0x00000168B5D23780> [label=Fare]
	<__main__.Node object at 0x00000168B5CAF0F0> -> <__main__.Node object at 0x00000168B5D23780> [label=1]
	<__main__.Node object at 0x00000168B5D23358> [label=Embarked]
	<__main__.Node object at 0x00000168B5D23780> -> <__main__.Node object at 0x00000168B5D23358> [label="upper class"]
	<__main__.Node object at 0x00000168B5D23A90> [label=Survived]
	<__main__.Node object at 0x00000168B5D23358> -> <__main__.Node object at 0x00000168B5D23A90> [label=S]
	<__main__.Node object at 0x00000168B5CDB240> [label=Death]
	<__main__.Node object at 0x00000168B5CAD320> -> <__main__.Node object at 0x00000168B5CDB240> [label=child]
	<__main__.Node object at 0x00000168B5CDBE48> [label=Survived]
	<__main__.Node object at 0x00000168B5CAD320> -> <__main__.Node object at 0x00000168B5CDBE48> [label=teen]
	<__main__.Node object at 0x00000168B5CFA908> [label=Parch]
	<__main__.Node object at 0x00000168B5C91780> -> <__main__.Node object at 0x00000168B5CFA908> [label=2]
	<__main__.Node object at 0x00000168B4C93470> [label=Embarked]
	<__main__.Node object at 0x00000168B5CFA908> -> <__main__.Node object at 0x00000168B4C93470> [label=0]
	<__main__.Node object at 0x00000168B5D23978> [label=Survived]
	<__main__.Node object at 0x00000168B4C93470> -> <__main__.Node object at 0x00000168B5D23978> [label=C]
	<__main__.Node object at 0x00000168B5D23048> [label=SibSp]
	<__main__.Node object at 0x00000168B4C93470> -> <__main__.Node object at 0x00000168B5D23048> [label=S]
	<__main__.Node object at 0x00000168B5D23B70> [label=Age]
	<__main__.Node object at 0x00000168B5D23048> -> <__main__.Node object at 0x00000168B5D23B70> [label=0]
	<__main__.Node object at 0x00000168B5D23C88> [label=Fare]
	<__main__.Node object at 0x00000168B5D23B70> -> <__main__.Node object at 0x00000168B5D23C88> [label=adults]
	<__main__.Node object at 0x00000168B5D23748> [label=Survived]
	<__main__.Node object at 0x00000168B5D23C88> -> <__main__.Node object at 0x00000168B5D23748> [label="middle class"]
	<__main__.Node object at 0x00000168B5D23EF0> [label=Survived]
	<__main__.Node object at 0x00000168B5D23B70> -> <__main__.Node object at 0x00000168B5D23EF0> [label=teen]
	<__main__.Node object at 0x00000168B5D23940> [label=Age]
	<__main__.Node object at 0x00000168B5D23048> -> <__main__.Node object at 0x00000168B5D23940> [label=1]
	<__main__.Node object at 0x00000168B5D23A20> [label=Fare]
	<__main__.Node object at 0x00000168B5D23940> -> <__main__.Node object at 0x00000168B5D23A20> [label=adults]
	<__main__.Node object at 0x00000168B5D23FD0> [label=Survived]
	<__main__.Node object at 0x00000168B5D23A20> -> <__main__.Node object at 0x00000168B5D23FD0> [label="middle class"]
	<__main__.Node object at 0x00000168B5D23828> [label=Survived]
	<__main__.Node object at 0x00000168B4C93470> -> <__main__.Node object at 0x00000168B5D23828> [label=Q]
	<__main__.Node object at 0x00000168B5D23C18> [label=SibSp]
	<__main__.Node object at 0x00000168B5CFA908> -> <__main__.Node object at 0x00000168B5D23C18> [label=1]
	<__main__.Node object at 0x00000168B5D232B0> [label=Survived]
	<__main__.Node object at 0x00000168B5D23C18> -> <__main__.Node object at 0x00000168B5D232B0> [label=0]
	<__main__.Node object at 0x00000168B5D234E0> [label=Age]
	<__main__.Node object at 0x00000168B5D23C18> -> <__main__.Node object at 0x00000168B5D234E0> [label=1]
	<__main__.Node object at 0x00000168B5D23E10> [label=Fare]
	<__main__.Node object at 0x00000168B5D234E0> -> <__main__.Node object at 0x00000168B5D23E10> [label=adults]
	<__main__.Node object at 0x00000168B5CAFCC0> [label=Embarked]
	<__main__.Node object at 0x00000168B5D23E10> -> <__main__.Node object at 0x00000168B5CAFCC0> [label="middle class"]
	<__main__.Node object at 0x00000168B5CDB198> [label=Survived]
	<__main__.Node object at 0x00000168B5CAFCC0> -> <__main__.Node object at 0x00000168B5CDB198> [label=S]
	<__main__.Node object at 0x00000168B5D23D68> [label=Survived]
	<__main__.Node object at 0x00000168B5D234E0> -> <__main__.Node object at 0x00000168B5D23D68> [label=child]
	<__main__.Node object at 0x00000168B5D23EB8> [label=Survived]
	<__main__.Node object at 0x00000168B5D23C18> -> <__main__.Node object at 0x00000168B5D23EB8> [label=2]
	<__main__.Node object at 0x00000168B5CADC18> [label=Survived]
	<__main__.Node object at 0x00000168B5CFA908> -> <__main__.Node object at 0x00000168B5CADC18> [label=2]
	<__main__.Node object at 0x00000168B5CAD0F0> [label=Survived]
	<__main__.Node object at 0x00000168B5CFA908> -> <__main__.Node object at 0x00000168B5CAD0F0> [label=3]
}
